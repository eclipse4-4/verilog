module syc_FIFO #(
    parameter DATA_WIDTH = 32,
    parameter DEPTH      = 8
)(
    input                       wr_en,
    input                       rd_en,
    input      [DATA_WIDTH-1:0] wr_data,
    input                       clk,
    input                       rstb,
    output reg [DATA_WIDTH-1:0] rd_data,
    output wire                 full,
    output wire                 empty
);

    // ????? ?? ???? localparam?? ???? ?? ? ??? ? ????.
    localparam ADDR_WIDTH = $clog2(DEPTH);
    localparam PTR_WIDTH  = ADDR_WIDTH + 1;

    // ?? ?? ??
    reg  [DATA_WIDTH-1:0] memory[DEPTH-1:0];
    reg  [PTR_WIDTH-1:0]  wr_ptr, rd_ptr;
    wire [DATA_WIDTH-1:0] rd_data_from_mem; // RAM ?? ?? ??? ?? wire

    // Full/Empty ?? (?? ?? ? ??? ??)
    assign full  = (wr_ptr[ADDR_WIDTH-1:0] == rd_ptr[ADDR_WIDTH-1:0]) &&
                   (wr_ptr[PTR_WIDTH-1]  != rd_ptr[PTR_WIDTH-1]);
    assign empty = (wr_ptr == rd_ptr);

    // === ??(Write) ?? - ??? always ???? ?? ===
    always @(posedge clk , negedge rstb) begin
        if (!rstb) begin
            wr_ptr <= 0;
        end else begin
            if (wr_en && !full) begin
                memory[wr_ptr[ADDR_WIDTH-1:0]] <= wr_data; // ???? ???
                wr_ptr <= wr_ptr + 1;
            end
        end
    end

    /* === ??(Read) ?? - ??? always ???? ?? ? ?? ?? ?? ===
    // 1. ????? ??? ???? (?? ?? ?? ?? ??)
     BRAM? ??? ??? ???: ??? ?? ???? ?? (???) MUX
     ?? ??????? read ??????? clk? ???, ??? clk?? ???? ???
     ????? ??? ???? ??? ???????? 1clk??? rd_data_from_mem? ?? ?? */
    assign rd_data_from_mem = memory[rd_ptr[ADDR_WIDTH-1:0]];

    // 2. ?? ?? ? ?? ??? ?????
    always @(posedge clk or negedge rstb) begin
        if (!rstb) begin
            rd_ptr  <= 0;
            rd_data <= 0;
        end else begin
            if (rd_en && !empty) begin
                rd_ptr  <= rd_ptr + 1;
                // ?? rd_ptr ??? ???? ???(rd_data_from_mem)? ?? ??? ???? ?? rd_data? ??
                rd_data <= rd_data_from_mem;
            end
        end
    end

endmodule

